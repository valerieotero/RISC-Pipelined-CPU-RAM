module ram256x32(output reg[31:0] DataOut, input Enable, ReadWrite, input [31:0] Address, input [31:0] DataIn)

endmodule 