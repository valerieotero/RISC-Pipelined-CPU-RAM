`include "mem.v"

module mem_tb;
endmodule